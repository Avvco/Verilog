module seven_segment_display(value, outSeg) ;
	input [3:0] value ;
	output [6:0] outSeg ;
	reg [6:0] outSeg ;
	always @(value)
	begin
		case(value)
			4'b0000: outSeg = 7'b1000000 ; // 0
			4'b0001: outSeg = 7'b1111001 ; // 1
			4'b0010: outSeg = 7'b0100100 ; // 2
			4'b0011: outSeg = 7'b0110000 ; // 3
			4'b0100: outSeg = 7'b0011001 ; // 4
			4'b0101: outSeg = 7'b0010010 ; // 5
			4'b0110: outSeg = 7'b0000010 ; // 6
			4'b0111: outSeg = 7'b1111000 ; // 7
			4'b1000: outSeg = 7'b0000000 ; // 8
			4'b1001: outSeg = 7'b0011000 ; // 9
			4'b1010: outSeg = 7'b0001000 ; // A
			4'b1011: outSeg = 7'b0000011 ; // b
			4'b1100: outSeg = 7'b1000110 ; // C
			4'b1101: outSeg = 7'b0100001 ; // d
			4'b1110: outSeg = 7'b0000110 ; // E
			4'b1111: outSeg = 7'b0001110 ; // F
		endcase
	end
endmodule